typedef uvm_sequencer #(empty_tx) empty_sequencer;




